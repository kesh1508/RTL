#work not_logic
#author keshave
#date 17-12-22
module not_logic (a_in, y_out);
input a_in;
output y_out;
assign y_out = ~a_in;
endmodule